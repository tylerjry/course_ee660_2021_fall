`timescale 1ns / 1ps

module lc4_divider(dividend_in, divisor_in, remainder_out, quotient_out);
   
   input [15:0] dividend_in, divisor_in;
   output [15:0] remainder_out, quotient_out;

   /*** YOUR CODE HERE ***/

endmodule


