`timescale 1ns / 1ps

module lc4_alu(insn, pc, r1data, r2data, out);
   
   input [15:0] insn, pc, r1data, r2data;
   output [15:0] out;
   
   /*** YOUR CODE HERE ***/

endmodule

